module transmitter(output logic tx);
initial
begin
tx<=1;
#1000000
$display("Frames: 0 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 2 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 3 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 4 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 5 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 6 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 7 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 8 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 9 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 10 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 11 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 12 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 13 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 14 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 15 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 16 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 17 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 18 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 19 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 20 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 21 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 22 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 23 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 24 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 25 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 26 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 27 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 28 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 29 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 30 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 31 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 32 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 33 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 34 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 35 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 36 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 37 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 38 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 39 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 40 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 41 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 42 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 43 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 44 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 45 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 46 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 47 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 48 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 49 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 50 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 51 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 52 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 53 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 54 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 55 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 56 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 57 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 58 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 59 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 60 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 61 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 62 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 63 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 64 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 65 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 66 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 67 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 68 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 69 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 70 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 71 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 72 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 73 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 74 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 75 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 76 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 77 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 78 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 79 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 80 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 81 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 82 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 83 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 84 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 85 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 86 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 87 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 88 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 89 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 90 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 91 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 92 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 93 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 94 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 95 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 96 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 97 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 98 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 99 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 100 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 101 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 102 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 103 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 104 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 105 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 106 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 107 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 108 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 109 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 110 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 111 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 112 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 113 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 114 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 115 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 116 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 117 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 118 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 119 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 120 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 121 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 122 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 123 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 124 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 125 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 126 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 127 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 128 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 129 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 130 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 131 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 132 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 133 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 134 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 135 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 136 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 137 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 138 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 139 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 140 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 141 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 142 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 143 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 144 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 145 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 146 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 147 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 148 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 149 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 150 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 151 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 152 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 153 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 154 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 155 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 156 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 157 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 158 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 159 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 160 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 161 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 162 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 163 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 164 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 165 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 166 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 167 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 168 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 169 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 170 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 171 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 172 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 173 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 174 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 175 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 176 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 177 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 178 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 179 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 180 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 181 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 182 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 183 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 184 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 185 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 186 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 187 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 188 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 189 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 190 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 191 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 192 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 193 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 194 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 195 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 196 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 197 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 198 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 199 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 200 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 201 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 202 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 203 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 204 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 205 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 206 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 207 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 208 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 209 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 210 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 211 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 212 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 213 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 214 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 215 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 216 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 217 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 218 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 219 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 220 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 221 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 222 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 223 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 224 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 225 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 226 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 227 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 228 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 229 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 230 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 231 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 232 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 233 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 234 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 235 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 236 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 237 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 238 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 239 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 240 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 241 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 242 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 243 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 244 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 245 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 246 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 247 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 248 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 249 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 250 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 251 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 252 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 253 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 254 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 255 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 256 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 257 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 258 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 259 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 260 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 261 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 262 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 263 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 264 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 265 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 266 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 267 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 268 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 269 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 270 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 271 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 272 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 273 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 274 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 275 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 276 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 277 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 278 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 279 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 280 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 281 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 282 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 283 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 284 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 285 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 286 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 287 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 288 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 289 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 290 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 291 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 292 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 293 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 294 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 295 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 296 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 297 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 298 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 299 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 300 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 301 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 302 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 303 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 304 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 305 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 306 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 307 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 308 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 309 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 310 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 311 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 312 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 313 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 314 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 315 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 316 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 317 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 318 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 319 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 320 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 321 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 322 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 323 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 324 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 325 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 326 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 327 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 328 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 329 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 330 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 331 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 332 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 333 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 334 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 335 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 336 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 337 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 338 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 339 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 340 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 341 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 342 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 343 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 344 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 345 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 346 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 347 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 348 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 349 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 350 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 351 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 352 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 353 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 354 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 355 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 356 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 357 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 358 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 359 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 360 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 361 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 362 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 363 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 364 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 365 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 366 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 367 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 368 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 369 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 370 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 371 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 372 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 373 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 374 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 375 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 376 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 377 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 378 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 379 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 380 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 381 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 382 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 383 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 384 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 385 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 386 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 387 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 388 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 389 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 390 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 391 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 392 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 393 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 394 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 395 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 396 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 397 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 398 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 399 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 400 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 401 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 402 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 403 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 404 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 405 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 406 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 407 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 408 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 409 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 410 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 411 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 412 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 413 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 414 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 415 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 416 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 417 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 418 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 419 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 420 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 421 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 422 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 423 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 424 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 425 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 426 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 427 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 428 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 429 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 430 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 431 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 432 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 433 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 434 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 435 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 436 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 437 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 438 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 439 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 440 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 441 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 442 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 443 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 444 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 445 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 446 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 447 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 448 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 449 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 450 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 451 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 452 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 453 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 454 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 455 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 456 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 457 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 458 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 459 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 460 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 461 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 462 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 463 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 464 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 465 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 466 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 467 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 468 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 469 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 470 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 471 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 472 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 473 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 474 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 475 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 476 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 477 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 478 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 479 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 480 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 481 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 482 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 483 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 484 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 485 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 486 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 487 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 488 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 489 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 490 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 491 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 492 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 493 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 494 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 495 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 496 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 497 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 498 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 499 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 500 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 501 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 502 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 503 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 504 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 505 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 506 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 507 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 508 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 509 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 510 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 511 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 512 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 513 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 514 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 515 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 516 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 517 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 518 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 519 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 520 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 521 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 522 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 523 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 524 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 525 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 526 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 527 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 528 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 529 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 530 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 531 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 532 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 533 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 534 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 535 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 536 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 537 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 538 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 539 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 540 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 541 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 542 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 543 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 544 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 545 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 546 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 547 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 548 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 549 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 550 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 551 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 552 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 553 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 554 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 555 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 556 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 557 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 558 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 559 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 560 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 561 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 562 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 563 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 564 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 565 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 566 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 567 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 568 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 569 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 570 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 571 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 572 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 573 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 574 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 575 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 576 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 577 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 578 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 579 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 580 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 581 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 582 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 583 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 584 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 585 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 586 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 587 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 588 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 589 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 590 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 591 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 592 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 593 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 594 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 595 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 596 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 597 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 598 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 599 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 600 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 601 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 602 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 603 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 604 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 605 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 606 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 607 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 608 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 609 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 610 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 611 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 612 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 613 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 614 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 615 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 616 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 617 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 618 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 619 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 620 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 621 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 622 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 623 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 624 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 625 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 626 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 627 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 628 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 629 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 630 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 631 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 632 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 633 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 634 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 635 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 636 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 637 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 638 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 639 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 640 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 641 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 642 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 643 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 644 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 645 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 646 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 647 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 648 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 649 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 650 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 651 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 652 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 653 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 654 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 655 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 656 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 657 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 658 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 659 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 660 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 661 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 662 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 663 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 664 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 665 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 666 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 667 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 668 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 669 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 670 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 671 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 672 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 673 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 674 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 675 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 676 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 677 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 678 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 679 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 680 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 681 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 682 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 683 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 684 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 685 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 686 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 687 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 688 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 689 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 690 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 691 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 692 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 693 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 694 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 695 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 696 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 697 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 698 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 699 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 700 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 701 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 702 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 703 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 704 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 705 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 706 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 707 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 708 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 709 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 710 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 711 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 712 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 713 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 714 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 715 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 716 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 717 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 718 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 719 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 720 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 721 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 722 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 723 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 724 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 725 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 726 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 727 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 728 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 729 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 730 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 731 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 732 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 733 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 734 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 735 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 736 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 737 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 738 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 739 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 740 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 741 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 742 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 743 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 744 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 745 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 746 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 747 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 748 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 749 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 750 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 751 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 752 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 753 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 754 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 755 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 756 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 757 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 758 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 759 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 760 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 761 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 762 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 763 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 764 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 765 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 766 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 767 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 768 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 769 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 770 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 771 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 772 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 773 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 774 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 775 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 776 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 777 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 778 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 779 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 780 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 781 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 782 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 783 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 784 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 785 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 786 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 787 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 788 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 789 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 790 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 791 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 792 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 793 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 794 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 795 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 796 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 797 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 798 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 799 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 800 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 801 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 802 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 803 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 804 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 805 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 806 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 807 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 808 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 809 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 810 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 811 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 812 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 813 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 814 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 815 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 816 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 817 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 818 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 819 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 820 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 821 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 822 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 823 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 824 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 825 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 826 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 827 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 828 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 829 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 830 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 831 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 832 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 833 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 834 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 835 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 836 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 837 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 838 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 839 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 840 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 841 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 842 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 843 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 844 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 845 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 846 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 847 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 848 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 849 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 850 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 851 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 852 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 853 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 854 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 855 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 856 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 857 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 858 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 859 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 860 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 861 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 862 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 863 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 864 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 865 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 866 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 867 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 868 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 869 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 870 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 871 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 872 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 873 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 874 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 875 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 876 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 877 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 878 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 879 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 880 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 881 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 882 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 883 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 884 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 885 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 886 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 887 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 888 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 889 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 890 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 891 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 892 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 893 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 894 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 895 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 896 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 897 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 898 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 899 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 900 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 901 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 902 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 903 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 904 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 905 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 906 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 907 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 908 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 909 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 910 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 911 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 912 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 913 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 914 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 915 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 916 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 917 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 918 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 919 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 920 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 921 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 922 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 923 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 924 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 925 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 926 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 927 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 928 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 929 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 930 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 931 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 932 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 933 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 934 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 935 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 936 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 937 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 938 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 939 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 940 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 941 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 942 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 943 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 944 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 945 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 946 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 947 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 948 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 949 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 950 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 951 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 952 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 953 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 954 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 955 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 956 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 957 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 958 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 959 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 960 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 961 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 962 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 963 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 964 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 965 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 966 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 967 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 968 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 969 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 970 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 971 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 972 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 973 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 974 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 975 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 976 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 977 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 978 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 979 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 980 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 981 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 982 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 983 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 984 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 985 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 986 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 987 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 988 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 989 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 990 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 991 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 992 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 993 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 994 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 995 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 996 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 997 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 998 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 999 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1000 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1001 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1002 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1003 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1004 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1005 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1006 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1007 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1008 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1009 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1010 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1011 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1012 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1013 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1014 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1015 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1016 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1017 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1018 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1019 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1020 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1021 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1022 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1023 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1024 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1025 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1026 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1027 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1028 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1029 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1030 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1031 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1032 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1033 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1034 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1035 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1036 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1037 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1038 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1039 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1040 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1041 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1042 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1043 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1044 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1045 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1046 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1047 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1048 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1049 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1050 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1051 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1052 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1053 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1054 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1055 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1056 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1057 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1058 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1059 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1060 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1061 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1062 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1063 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1064 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1065 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1066 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1067 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1068 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1069 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1070 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1071 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1072 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1073 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1074 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1075 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1076 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1077 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1078 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1079 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1080 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1081 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1082 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1083 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1084 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1085 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1086 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1087 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1088 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1089 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1090 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1091 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1092 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1093 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1094 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1095 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1096 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1097 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1098 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1099 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1100 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1101 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1102 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1103 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1104 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1105 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1106 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1107 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1108 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1109 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1110 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1111 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1112 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1113 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1114 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1115 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1116 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1117 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1118 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1119 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1120 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1121 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1122 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1123 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1124 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1125 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1126 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1127 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1128 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1129 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1130 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1131 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1132 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1133 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1134 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1135 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1136 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1137 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1138 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1139 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1140 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1141 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1142 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1143 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1144 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1145 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1146 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1147 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1148 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1149 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1150 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1151 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1152 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1153 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1154 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1155 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1156 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1157 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1158 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1159 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1160 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1161 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1162 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1163 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1164 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1165 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1166 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1167 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1168 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1169 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1170 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1171 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1172 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1173 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1174 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1175 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1176 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1177 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1178 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1179 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1180 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1181 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1182 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1183 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1184 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1185 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1186 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1187 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1188 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1189 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1190 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1191 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1192 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1193 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1194 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1195 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1196 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1197 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1198 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1199 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1200 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1201 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1202 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1203 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1204 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1205 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1206 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1207 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1208 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1209 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1210 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1211 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1212 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1213 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1214 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1215 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1216 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1217 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1218 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1219 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1220 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1221 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1222 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1223 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1224 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1225 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1226 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1227 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1228 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1229 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1230 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1231 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1232 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1233 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1234 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1235 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1236 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1237 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1238 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1239 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1240 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1241 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1242 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1243 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1244 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1245 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1246 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1247 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1248 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1249 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1250 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1251 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1252 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1253 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1254 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1255 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1256 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1257 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1258 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1259 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1260 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1261 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1262 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1263 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1264 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1265 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1266 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1267 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1268 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1269 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1270 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1271 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1272 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1273 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1274 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1275 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1276 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1277 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1278 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1279 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1280 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1281 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1282 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1283 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1284 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1285 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1286 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1287 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1288 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1289 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1290 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1291 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1292 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1293 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1294 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1295 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1296 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1297 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1298 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1299 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1300 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1301 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1302 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1303 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1304 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1305 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1306 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1307 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1308 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1309 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1310 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1311 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1312 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1313 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1314 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1315 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1316 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1317 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1318 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1319 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1320 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1321 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1322 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1323 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1324 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1325 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1326 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1327 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1328 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1329 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1330 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1331 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1332 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1333 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1334 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1335 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1336 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1337 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1338 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1339 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1340 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1341 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1342 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1343 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1344 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1345 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1346 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1347 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1348 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1349 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1350 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1351 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1352 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1353 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1354 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1355 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1356 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1357 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1358 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1359 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1360 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1361 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1362 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1363 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1364 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1365 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1366 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1367 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1368 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1369 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1370 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1371 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1372 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1373 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1374 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1375 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1376 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1377 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1378 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1379 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1380 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1381 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1382 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1383 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1384 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1385 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1386 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1387 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1388 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1389 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1390 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1391 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1392 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1393 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1394 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1395 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1396 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1397 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1398 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1399 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1400 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1401 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1402 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1403 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1404 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1405 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1406 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1407 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1408 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1409 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1410 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1411 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1412 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1413 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1414 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1415 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1416 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1417 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1418 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1419 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1420 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1421 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1422 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1423 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1424 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1425 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1426 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1427 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1428 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1429 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1430 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1431 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1432 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1433 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1434 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1435 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1436 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1437 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1438 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1439 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1440 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1441 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1442 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1443 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1444 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1445 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1446 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1447 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
$display("Frames: 1448 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1449 / 1450");
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 0;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
#200 tx <= 1;
$display("Frames: 1450 / 1450");
#200 tx<=1;
#1000000 $finish;
end
endmodule